module bb_iocell (
    inout vdd,
    inout vss,
    inout vddio,
    inout vssio,
    inout poc
);

endmodule