(* blackbox *) 
module IOPAD (
    input A,
    input EN,
    output Y,
    inout PAD
);

endmodule